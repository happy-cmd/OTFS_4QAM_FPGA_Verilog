`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/11/15 16:55:36
// Design Name: 
// Module Name: OTFSTx_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//--------------------------------------------------------------------------------------------
//
// Generated by X-HDL VHDL Translator - Version 2.0.0 Feb. 1, 2011
// ?? 10? 31 2024 11:14:47
//
//      Input file      : 
//      Component name  : otfstx
//      Author          : 
//      Company         : 
//
//      Description     : 
//
//
//--------------------------------------------------------------------------------------------


module OTFSTx_32(Clk, SRst, Start, DataValid, DataIn, ModDataOutValid, FrameBeginnigIndicator, FrameNum, DataNum, ModDataOutRe, ModDataOutIm, OTFSTxDataValid, OTFSTxDataRe, OTFSTxDataIm);
   input         Clk;
   input         SRst;
   input         Start;
   
   input         DataValid;
   input         DataIn;
   
   output        ModDataOutValid;
   output        FrameBeginnigIndicator;
   output [7:0]  FrameNum;
   output [7:0]  DataNum;
   output [11:0] ModDataOutRe;
   output [11:0] ModDataOutIm;
   
   output        OTFSTxDataValid;
   output [15:0] OTFSTxDataRe;
   output [15:0] OTFSTxDataIm;
   
   
   wire [11:0]   ModDataOutReReg;
   wire [11:0]   ModDataOutImReg;
   wire          ModDataOutValidReg;
   wire [1:0]   QAMData_instruct;
   
   assign ModDataOutRe = ModDataOutReReg;
   assign ModDataOutIm = ModDataOutImReg;
   assign ModDataOutValid = ModDataOutValidReg;
   
   QAMModulator_32QAM U1(
   .Clk(Clk), 
   .SRst(SRst), 
   .Start(Start), 
   .DataValidIn(DataValid), 
   .Data(DataIn), 
   .ModDataOutValid(ModDataOutValidReg), 
   .FrameBeginnigIndicator(FrameBeginnigIndicator), 
   .FrameNum(FrameNum), 
   .DataNum(DataNum), 
   .ModDataOutRe(ModDataOutReReg), 
   .ModDataOutIm(ModDataOutImReg)
   );
   
   
   OTFSModulator U2(
   .Clk(Clk), 
   .Srst(SRst), 
   .Start(Start), 
   .QAMDataValid(ModDataOutValidReg), 
   .QAMDataRe(ModDataOutReReg), 
   .QAMDataIm(ModDataOutImReg), 
   .OTFSTxDataValid(OTFSTxDataValid), 
   .OTFSTxDataRe(OTFSTxDataRe), 
   .OTFSTxDataIm(OTFSTxDataIm)
   );
   
endmodule
