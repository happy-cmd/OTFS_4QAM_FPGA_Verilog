`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/11/15 16:38:16
// Design Name: 
// Module Name: TopModule_Verilog
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//--------------------------------------------------------------------------------------------
//
// Generated by X-HDL VHDL Translator - Version 2.0.0 Feb. 1, 2011
// ?? 10? 31 2024 11:14:30
//
//      Input file      : 
//      Component name  : topmodule
//      Author          : 
//      Company         : 
//
//      Description     : 
//
//
//--------------------------------------------------------------------------------------------


module TopModule_Verilog (
    Clk,
    SRst,
    Start,
    ModulationOrder,
    QAMModDataOutValid,
    QAMFrameBeginnigIndicator,
    QAMFrameNum,
    QAMDataNum,
    QAMModDataOutRe,
    QAMModDataOutIm,
    OTFSTxDataValid,
    OTFSTxDataRe,
    OTFSTxDataIm,
    OTFSRxDemodValid,
    OTFSRxDemodRe,
    OTFSRxDemodIm,
    QAMDemodDataValid,
    QAMDemodData
);
  input Clk;
  input SRst;
  input Start;
  input [2:0] ModulationOrder;

  output QAMModDataOutValid;
  output QAMFrameBeginnigIndicator;
  output [7:0] QAMFrameNum;
  output [7:0] QAMDataNum;
  output [11:0] QAMModDataOutRe;
  output [11:0] QAMModDataOutIm;

  output OTFSTxDataValid;
  output [15:0] OTFSTxDataRe;
  output [15:0] OTFSTxDataIm;

  output OTFSRxDemodValid;
  output [23:0] OTFSRxDemodRe;
  output [23:0] OTFSRxDemodIm;

  output QAMDemodDataValid;
  output [4:0] QAMDemodData;


  wire        RandomBitValid;
  wire        RandomBit;

  wire        ModDataOutValidReg;
  wire        FrameBeginnigIndicatorReg;
  wire [ 7:0] FrameNumReg;
  wire [ 7:0] DataNumReg;
  wire [11:0] ModDataOutReReg;
  wire [11:0] ModDataOutImReg;
  wire        OTFSDataValidReg;
  wire [15:0] OTFSDataReReg;
  wire [15:0] OTFSDataImReg;


  RandomBitGenerator U0 (
      .Clk(Clk),
      .SRst(SRst),
      .Start(Start),
      .ModulationOrder(ModulationOrder),
      .RandomBitValid(RandomBitValid),
      .RandomBit(RandomBit)
  );
  
       integer handle1;
      initial
      begin
       handle1 =  $fopen("../../../../../sim_result/RandomBit_Gene_32QAM.txt");
      end
      always@(posedge Clk)
      begin
        if(RandomBitValid)
          begin
            $fdisplay(handle1,"%d",RandomBit);
          end
      end

  assign QAMModDataOutValid = ModDataOutValidReg;
  assign QAMFrameBeginnigIndicator = FrameBeginnigIndicatorReg;
  assign QAMFrameNum = FrameNumReg;
  assign QAMDataNum = DataNumReg;
  assign QAMModDataOutRe = ModDataOutReReg;
  assign QAMModDataOutIm = ModDataOutImReg;

  assign OTFSTxDataValid = OTFSDataValidReg;
  assign OTFSTxDataRe = OTFSDataReReg;
  assign OTFSTxDataIm = OTFSDataImReg;


  OTFSTx_32 U1 (
      .Clk(Clk),
      .SRst(SRst),
      .Start(Start),
      .DataValid(RandomBitValid),
      .DataIn(RandomBit),
      .ModDataOutValid(ModDataOutValidReg),
      .FrameBeginnigIndicator(FrameBeginnigIndicatorReg),
      .FrameNum(FrameNumReg),
      .DataNum(DataNumReg),
      .ModDataOutRe(ModDataOutReReg),
      .ModDataOutIm(ModDataOutImReg),
      .OTFSTxDataValid(OTFSDataValidReg),
      .OTFSTxDataRe(OTFSDataReReg),
      .OTFSTxDataIm(OTFSDataImReg)
  );
  
       integer handle2,handle3;
      initial
      begin
       handle2 =  $fopen("../../../../../sim_result/QAMModDataOutRe_32QAM.txt");
       handle3 =  $fopen("../../../../../sim_result/QAMModDataOutIm_32QAM.txt");
      end
      always@(posedge Clk)
      begin
        if(QAMModDataOutValid)
          begin
            $fdisplay(handle2,"%d",$signed(QAMModDataOutRe));
            $fdisplay(handle3,"%d",$signed(QAMModDataOutIm));
          end
      end
      
      integer handle4;
      initial
      begin
       handle4 =  $fopen("../../../../../sim_result/OTFSModResult_32QAM.txt");
      end
      always@(posedge Clk)
      begin
        if(OTFSTxDataValid)
          begin
            $fdisplay(handle4,"%d,%d", $signed(OTFSTxDataRe), $signed(OTFSTxDataIm));
          end
      end
  OTFSRx_32 U2 (
      .Clk(Clk),
      .Srst(SRst),
      .Start(Start),
      .RecSigDataValid(OTFSDataValidReg),
      .RecSigRe(OTFSDataReReg),
      .RecSigIm(OTFSDataImReg),
      .OTFSRxDemodValid(OTFSRxDemodValid),
      .OTFSRxDemodRe(OTFSRxDemodRe),
      .OTFSRxDemodIm(OTFSRxDemodIm),
      .QAMDemodDataValid(QAMDemodDataValid),
      .QAMDemodData(QAMDemodData)
  );
 integer handle5;
  initial
  begin
   handle5 =  $fopen("../../../../../sim_result/OTFSDeModResult_32QAM.txt");
  end
  always@(posedge Clk)
  begin
    if(OTFSRxDemodValid)
      begin
        $fdisplay(handle5,"%d,%d", $signed(OTFSRxDemodRe), $signed(OTFSRxDemodIm));
      end
  end
  
integer handle6,handle7;
 initial
 begin
  handle6 =  $fopen("../../../../../sim_result/QAMDeModDataOut_32QAM.txt");
 end
 always@(posedge Clk)
 begin
   if(QAMDemodDataValid)
     begin
       $fdisplay(handle6,"%d",$unsigned(QAMDemodData));
     end
 end
endmodule
